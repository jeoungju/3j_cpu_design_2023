module p_d_MW(
    port_list
);
    
endmodule