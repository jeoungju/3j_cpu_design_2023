module p_d_EM(
    port_list
);
    
endmodule