//`timescale 1ns/1ps

`include "opcode.vh"
`include "mem_path.vh"

// This testbench tests if the cpu module can decode and execute
// all the instructions specified in the spec (RV32I -- including CSRRW and CSRRWI).
// Some tests for data hazards and control hazards are also included.

// How does the testbench work?
// For each test, the testbench initializes IMem with one or several instructions
// (encoded in binary format as specified in the spec) for testing.
// RegFile and DMem are also initialized with some data.
// Then, the clock is advanced until the cpu module gives correct result
// in the RegFile or DMem. If no correct result is returned after a "timeout" cycle,
// the testbench will be terminated (or failed)

// This setting is different from other testbenches, in which the BIOSMem or IMem is initialized
// with a hex file generated by compiling the assembly/C code of the corresponding
// test software (the hex file contains the binary encoding of the instructions and data
// of the program). Here, we manually generate the instructions and data.

// Don't just run the testbench, look at the tests, see what they do.
// The testbench is intended to provide you some examples to get started.
// Feel free to make your own change.
// Note that the testbench is by no means exhaustive.
// You should add your own tests if there are cases you think the testbench
// does not cover.

module cpu_tb();
  reg clk, rst;
  parameter CPU_CLOCK_PERIOD = 20;
  parameter CPU_CLOCK_FREQ   = 1_000_000_000 / CPU_CLOCK_PERIOD;

  initial clk = 0;
  always #(CPU_CLOCK_PERIOD/2) clk = ~clk;
  wire [31:0] csr;

  // Init PC with 32'h1000_0000 -- address space of IMem
  // When PC is in IMem's address space, IMem is read-only
  // DMem can be R/W as long as the addr bits [31:28] is 4'b00x1
  // cpu # (
  //   .CPU_CLOCK_FREQ(CPU_CLOCK_FREQ),
  //   .RESET_PC(32'h1000_0000)
  // ) CPU (
  //   .clk(clk),
  //   .rst(rst),
  //   .serial_in(1'b1),
  //   .serial_out()
  // );

  // instantiate device to be tested
  // Reset: Low Active
  top #(
      .RESET_PC(32'h1000_0000),
      .MIF_HEX("")
  ) CPU (
      .clk    (clk),
      .n_rst  (~rst),
        .PC        (),
        .Instr     (),
      .WriteData (),
      .DataAdr   (),
      .MemWrite  ()
    );


  wire [31:0] timeout_cycle = 25; //10

  // Reset IMem, DMem, and RegFile before running new test
  task reset;
    integer i;
    begin
      for (i = 0; i < `RF_PATH.DEPTH; i = i + 1) begin
        `RF_PATH.mem[i] = 0;
      end
      for (i = 0; i < `DMEM_PATH.DEPTH; i = i + 1) begin
        `DMEM_PATH.mem[i] = 0;
      end
      for (i = 0; i < `IMEM_PATH.DEPTH; i = i + 1) begin
        `IMEM_PATH.mem[i] = 0;
      end
    end
  endtask

  task reset_cpu; 
      begin
    repeat (3) begin
      @(negedge clk);
      rst = 1;
    end
    @(negedge clk);
    rst = 0;
end
  endtask

  task init_rf;
    integer i;
    begin
      for (i = 1; i < `RF_PATH.DEPTH; i = i + 1) begin
        `RF_PATH.mem[i] = 100 * i + 1;
      end
    end
  endtask

  reg [31:0] cycle;
  reg done;
  reg [31:0]  current_test_id = 0;
  reg [255:0] current_test_type;
  reg [31:0]  current_output;
  reg [31:0]  current_result;
  reg all_tests_passed = 0;


  // Check for timeout
  // If a test does not return correct value in a given timeout cycle,
  // we terminate the testbench
  initial begin
    while (all_tests_passed === 0) begin
      @(posedge clk);
      if (cycle === timeout_cycle) begin
        $display("[Failed] Timeout at [%d] test %s, expected_result = %h, got = %h",
                current_test_id, current_test_type, current_result, current_output);
        $finish();
      end
    end
  end

  always @(posedge clk) begin
    if (done === 0)
      cycle <= cycle + 1;
    else
      cycle <= 0;
  end

  // Check result of RegFile
  // If the write_back (destination) register has correct value (matches "result"), test passed
  // This is used to test instructions that update RegFile
  task check_result_rf;
    input [31:0]  rf_wa;
    input [31:0]  result;
    input [255:0] test_type;
    begin
      done = 0;
      current_test_id   = current_test_id + 1;
      current_test_type = test_type;
      current_result    = result;
      while (`RF_PATH.mem[rf_wa] !== result) begin
        current_output = `RF_PATH.mem[rf_wa];
        @(posedge clk);
      end
      cycle = 0;
      done = 1;
      $display("[%d] Test %s passed!", current_test_id, test_type);
    end
  endtask

  // Check result of DMem
  // If the memory location of DMem has correct value (matches "result"), test passed
  // This is used to test store instructions
  task check_result_dmem;
    input [31:0]  addr;
    input [31:0]  result;
    input [255:0] test_type;
    begin
      done = 0;
      current_test_id   = current_test_id + 1;
      current_test_type = test_type;
      current_result    = result;
      while (`DMEM_PATH.mem[addr] !== result) begin
        current_output = `DMEM_PATH.mem[addr];
        @(posedge clk);
      end
      cycle = 0;
      done = 1;
      $display("[%d] Test %s passed!", current_test_id, test_type);
    end
  endtask

  integer i;

  reg [31:0] num_cycles = 0;
  reg [31:0] num_insts  = 0;
  reg [4:0]  RD, RS1, RS2, RS3;
  reg [31:0] RD1, RD2, RD3;
  reg [4:0]  SHAMT;
  reg [31:0] IMM, IMM0, IMM1, IMM2, IMM3;
  reg [14:0] INST_ADDR;
  reg [14:0] DATA_ADDR;
  reg [14:0] DATA_ADDR0, DATA_ADDR1, DATA_ADDR2, DATA_ADDR3;
  reg [14:0] DATA_ADDR4, DATA_ADDR5, DATA_ADDR6, DATA_ADDR7;
  reg [14:0] DATA_ADDR8, DATA_ADDR9;

  reg [31:0] JUMP_ADDR, AFTER_ADDR;

  reg [31:0]  BR_TAKEN_OP1  [5:0];
  reg [31:0]  BR_TAKEN_OP2  [5:0];
  reg [31:0]  BR_NTAKEN_OP1 [5:0];
  reg [31:0]  BR_NTAKEN_OP2 [5:0];
  reg [2:0]   BR_TYPE       [5:0];
  reg [255:0] BR_NAME_TK1   [5:0];
  reg [255:0] BR_NAME_TK2   [5:0];
  reg [255:0] BR_NAME_NTK   [5:0];

  initial begin
    `ifndef IVERILOG
        $vcdpluson;
    `endif
    `ifdef IVERILOG
        $dumpfile("cpu_tb.fst");
        $dumpvars(0, cpu_tb);
    `endif
    `ifdef FSDB
        $fsdbDumpfile("wave.fsdb");
        $fsdbDumpvars(0);
    `endif

    #0;
    rst = 0;

    // Reset the CPU
    rst = 1;
    // Hold reset for a while
    repeat (10) @(posedge clk);

    @(negedge clk);
    rst = 0;

/*
if (1) begin
   // Test CSR Insts -----------------------------------------------------
   // - CSRRW, CSRRWI
  reset();

  `RF_PATH.mem[1] = 100;
  IMM       = 5'd16;
  INST_ADDR = 14'h0000;

  `IMEM_PATH.mem[INST_ADDR + 0] = {12'h51e, 5'd1,     3'b001, 5'd0, `OPC_CSR};
  `IMEM_PATH.mem[INST_ADDR + 1] = {12'h51e, IMM[4:0], 3'b101, 5'd0, `OPC_CSR};

  reset_cpu();

  current_test_id = current_test_id + 1;
  current_test_type = "CSRRW Test";
  done = 0;
  while (`CSR_PATH !== `RF_PATH.mem[1])
    @(posedge clk);
  done = 1;

  $display("[%d] Test CSRRW passed!", current_test_id);

  current_test_id = current_test_id + 1;
  current_test_type = "CSRRWI Test";
  done = 0;
  wait (`CSR_PATH === IMM);
  done = 1;

  $display("[%d] Test CSRRWI passed!", current_test_id);
end
*/

    // Your own Testbench
    // Add two testvector: each instruction
    // Add Instruction : -10 + 20 = 10

    // Test case 1
    reset();

    // We can also use $random to generate random values for testing
    /*
    RS1 = 1; RD1 = -10;
    RS2 = 2; RD2 =  20;
    RD  = 4;
    `RF_PATH.mem[RS1] = RD1;
    `RF_PATH.mem[RS2] = RD2;
    SHAMT           = 5'd20;
    INST_ADDR       = 14'h0000;

    `IMEM_PATH.mem[INST_ADDR + 0]  = {`FNC7_0, RS2,   RS1, `FNC_ADD_SUB, RD,  `OPC_ARI_RTYPE};

    reset_cpu();

    check_result_rf(RD,  32'h0000000a, "R-Type ADD");
    $display("[INFO: My CPU]Add Instruction Pass");
    */

    // Test case 2: Midterm Project
    //-------------------Start !!---------------------------
    if (1) begin
    // Test R-Type Insts --------------------------------------------------
    // - ADD, SUB, SLL, SLT, SLTU, SRL, SRA
    reset();

    // We can also use $random to generate random values for testing
    RS1 = 1; RD1 =  32'h7fff_ffff;
    RS2 = 2; RD2 =  32'h0000_0001;
    RS3 = 3; RD3 =  32'h8fff_ffff;
    RD  = 5;
    `RF_PATH.mem[RS1] = RD1; //x1 data
    `RF_PATH.mem[RS2] = RD2; //x2 data
    `RF_PATH.mem[RS3] = RD3; //x3 data
    INST_ADDR       = 14'h0000;

    `IMEM_PATH.mem[INST_ADDR + 0]  = {`FNC7_0, RS2,   RS1, `FNC_ADD_SUB, RD,  `OPC_ARI_RTYPE};
    //ADD x5, x1, x2 => x5 = 0x7fff_ffff + 0x0000_0001 = 32'h8000_0000 sign bit change overflow 
    `IMEM_PATH.mem[INST_ADDR + 1]  = {`FNC7_1, RS2,   RS1, `FNC_ADD_SUB, 5'd6,  `OPC_ARI_RTYPE};
    //SUB x6, x1, x2 => x6 = 0x7fff_ffff - 0x0000_0001 = 32'h7fff_fffe
    `IMEM_PATH.mem[INST_ADDR + 2]  = {`FNC7_0, RS2,   RS1, `FNC_SLL,     5'd7,  `OPC_ARI_RTYPE};
    //SLL x7, x1, x2 => x7 = x1(0x7fff_ffff) << x2[4:0](1) = 32'hffff_fffe
    `IMEM_PATH.mem[INST_ADDR + 3]  = {`FNC7_0, RS2,   RS3, `FNC_SLT,     5'd8,  `OPC_ARI_RTYPE};
    //SLT x8, x3, x2 => x3 -x2 < 0 ? 32'h1 : 32'h0 , x8 = 32'h1   // signed
    `IMEM_PATH.mem[INST_ADDR + 4]  = {`FNC7_0, RS2,   RS3, `FNC_SLTU,    5'd9,  `OPC_ARI_RTYPE};
    //SLTU x9, x3, x2 => x3 -x2 < 0 ? 32'h1 : 32'h0 , x9 = 32'h0 // unsigned
    `IMEM_PATH.mem[INST_ADDR + 5]  = {`FNC7_0, RS2,   RS3, `FNC_SRL_SRA, 5'd10, `OPC_ARI_RTYPE};
    //SRL x10, x3, x2 => x10 = x3(0x8fff_ffff) >> x2[4:0](1) = 32'h47ff_ffff //zero extension
    `IMEM_PATH.mem[INST_ADDR + 6]  = {`FNC7_1, RS2,   RS3, `FNC_SRL_SRA, 5'd11, `OPC_ARI_RTYPE};
    //SRA x11, x3, x2 => x11 = x3(0x8fff_ffff) >>> x2[4:0](1) = 32'hc7ff_ffff // sign extension

    reset_cpu();

    check_result_rf(RD,  32'h8000_0000, "R-Type ADD");
    check_result_rf(5'd6,  32'h7fff_fffe, "R-Type SUB");
    check_result_rf(5'd7,  32'hffff_fffe, "R-Type SLL");
    check_result_rf(5'd8,  32'h1,        "R-Type SLT");
    check_result_rf(5'd9,  32'h0,        "R-Type SLTU");
    check_result_rf(5'd10, 32'h47ff_ffff, "R-Type SRL");
    check_result_rf(5'd11, 32'hc7ff_ffff, "R-Type SRA");

end

if (1) begin
    // Test R-Type Insts --------------------------------------------------
    // - XOR, OR, AND

    reset();

    // We can also use $random to generate random values for testing
    RS1 = 1; RD1 = 32'hf0f0_a0a0;
    RS2 = 2; RD2 =  32'h0f0f_f0f0;
    RD  = 3;
    `RF_PATH.mem[RS1] = RD1;
    `RF_PATH.mem[RS2] = RD2;
    SHAMT           = 5'd20;
    INST_ADDR       = 14'h0000;

    `IMEM_PATH.mem[INST_ADDR + 0]  = {`FNC7_0, RS2,   RS1, `FNC_XOR,     5'd8,  `OPC_ARI_RTYPE};
    //XOR x8, x1, x2 => x8 = x1 ^ x2 = 0xf0f0_a0a0 ^ 0x0f0f_f0f0 = 0xffff_5050
    `IMEM_PATH.mem[INST_ADDR + 1]  = {`FNC7_0, RS2,   RS1, `FNC_OR,      5'd9,  `OPC_ARI_RTYPE};
    //OR x9, x1, x2 => x9 = x1 | x2 = 0xf0f0_a0a0 | 0x0f0f_f0f0 = 0xffff_f0f0
    `IMEM_PATH.mem[INST_ADDR + 2]  = {`FNC7_0, RS2,   RS1, `FNC_AND,     5'd10, `OPC_ARI_RTYPE};
    //AND x10, x1, x2 => x10 = x1 & x2 =  0xf0f0_a0a0 & 0x0f0f_f0f0 = 0x0000_a0a0


    reset_cpu();

    check_result_rf(5'd8,  32'hffff_5050, "R-Type XOR");
    check_result_rf(5'd9,  32'hffff_f0f0, "R-Type OR");
    check_result_rf(5'd10, 32'h0000_a0a0, "R-Type AND");

end

if (1) begin
    // Test I-Type Insts --------------------------------------------------
    // - ADDI, SLTI, SLTUI, XORI, ORI, ANDI
    // - LW, LH, LB, LHU, LBU
    // - JALR

    // Test I-type arithmetic instructions
    reset();

    RS1 = 1; RD1 = 32'hffff_ffe2; //-30  unsigned big data
    `RF_PATH.mem[RS1] = RD1;
    IMM             = 32'h0000_0014;  //20
    INST_ADDR       = 14'h0000;
    SHAMT           = 5'd16;

    `IMEM_PATH.mem[INST_ADDR + 0] = {IMM[11:0], RS1, `FNC_ADD_SUB, 5'd3, `OPC_ARI_ITYPE};
    //ADDI x3, x1, 20 => x3 = x1(-30) + 20 = -10(0xffff_fff6)
    `IMEM_PATH.mem[INST_ADDR + 1] = {IMM[11:0], RS1, `FNC_SLT,     5'd4, `OPC_ARI_ITYPE};
    //SLTI x4, x1, 20 => x1 -20 < 0 ? 1 : 0  //signed
    `IMEM_PATH.mem[INST_ADDR + 2] = {IMM[11:0], RS1, `FNC_SLTU,    5'd5, `OPC_ARI_ITYPE};
    //SLTUI x5, x1, 20 => x1 - 20 < 0 ? 1 : 0  //unsigned
    `IMEM_PATH.mem[INST_ADDR + 3] = {IMM[11:0], RS1, `FNC_XOR,     5'd6, `OPC_ARI_ITYPE};
    //XORI x6, x1, 20 => x6 = x1 ^ 20 = 0xffff_ffe2 ^ 0x0000_0014 = 0xffff_fff6
    `IMEM_PATH.mem[INST_ADDR + 4] = {IMM[11:0], RS1, `FNC_OR,      5'd7, `OPC_ARI_ITYPE};
    //ORI x7, x1, 20 => x7 = x1 | 20 = 0xffff_ffe2 | 0x0000_0014 = 0xffff_fff6
    `IMEM_PATH.mem[INST_ADDR + 5] = {IMM[11:0], RS1, `FNC_AND,     5'd8, `OPC_ARI_ITYPE};
    //ANDI x8, x1, 20 => x8 = x1 & 20 = 0xffff_ffe2 & 0x0000_0014 = 0x0000_0000 
    `IMEM_PATH.mem[INST_ADDR + 6] = {`FNC7_0, SHAMT, RS1, `FNC_SLL,     5'd9, `OPC_ARI_ITYPE};
    //SLLI x9, x1, 16 => x9 = x1 << 16 = 0xffff_ffe2 << 16 = 0xffe2_0000
    `IMEM_PATH.mem[INST_ADDR + 7] = {`FNC7_0, SHAMT, RS1, `FNC_SRL_SRA, 5'd10, `OPC_ARI_ITYPE};
    //SRLI x10, x1, 16 => x10 =  x1 >> 16 = 0xffff_ffe2 >> 16 = 0x0000_ffff //zero extension
    `IMEM_PATH.mem[INST_ADDR + 8] = {`FNC7_1, SHAMT, RS1, `FNC_SRL_SRA, 5'd11, `OPC_ARI_ITYPE};
    //SRAI x11, x1, 16 => x11 =  x1 >>> 16 = 0xffff_ffe2 >>> 16 = 0xffff_ffff //sign extension

    reset_cpu();

    check_result_rf(5'd3,  32'hffff_fff6, "I-Type ADDI");
    check_result_rf(5'd4,  32'h00000001, "I-Type SLTI");
    check_result_rf(5'd5,  32'h00000000, "I-Type SLTUI");
    check_result_rf(5'd6,  32'hffff_fff6, "I-Type XORI");
    check_result_rf(5'd7,  32'hffff_fff6, "I-Type ORI");
    check_result_rf(5'd8,  32'h0000_0000, "I-Type ANDI");
    check_result_rf(5'd9, 32'hffe2_0000, "I-Type SLLI"); //shamt = 16  0x10
    check_result_rf(5'd10, 32'h0000_ffff, "I-Type SRLI");
    check_result_rf(5'd11, 32'hffff_ffff, "I-Type SRAI");
end

if (1) begin
    // Test I-type load instructions
    reset();

    `RF_PATH.mem[1] = 32'h3000_0100; //x1 = 0x3000_0100, Data memory addr
    IMM0            = 32'h0000_0000; //Lasr Addr [1:0]
    IMM1            = 32'h0000_0001;
    IMM2            = 32'h0000_0002;
    IMM3            = 32'h0000_0003;
    INST_ADDR       = 14'h0000;
    DATA_ADDR       = (`RF_PATH.mem[1] + IMM0[11:0]) >> 2; 

    `IMEM_PATH.mem[INST_ADDR + 0] = {IMM0[11:0], 5'd1, `FNC_LW,  5'd2,  `OPC_LOAD};
    //LW x2, 0[x1] => x2 = mem[x1 + 0x000] = 32'hface_cafe
    `IMEM_PATH.mem[INST_ADDR + 1] = {IMM0[11:0], 5'd1, `FNC_LH,  5'd3,  `OPC_LOAD};
    //LH x3, 0[x1] => x3 = mem[x1 + 0x000] = 32'hffff_cafe
    `IMEM_PATH.mem[INST_ADDR + 2] = {IMM2[11:0], 5'd1, `FNC_LH,  5'd4,  `OPC_LOAD};
    //LH x4, 2[x1] => x4 = mem[x1 + 0x002] = 32'hffff_face
    `IMEM_PATH.mem[INST_ADDR + 3] = {IMM0[11:0], 5'd1, `FNC_LB,  5'd5,  `OPC_LOAD};
    //LB x5, 0[x1] => x5 = mem[x1 + 0x000] = 32'hffff_fffe
    `IMEM_PATH.mem[INST_ADDR + 4] = {IMM1[11:0], 5'd1, `FNC_LB,  5'd6,  `OPC_LOAD};
    //LB x6, 1[x1] => x6 = mem[x1 + 0x001] = 32'hffff_ffca
    `IMEM_PATH.mem[INST_ADDR + 5] = {IMM2[11:0], 5'd1, `FNC_LB,  5'd7,  `OPC_LOAD};
    //LB x7, 2[x1] => x7 = mem[x1 + 0x002] = 32'hffff_ffce
    `IMEM_PATH.mem[INST_ADDR + 6] = {IMM3[11:0], 5'd1, `FNC_LB,  5'd8, `OPC_LOAD};
    //LB x8, 3[x1] => x8 = mem[x1 + 0x003] = 32'hffff_fffa
    `IMEM_PATH.mem[INST_ADDR + 7] = {IMM0[11:0], 5'd1, `FNC_LHU, 5'd9, `OPC_LOAD};
    //LHU x9, 0[x1] => x9 = mem[x1 + 0x000] = 32'h0000_cafe
    `IMEM_PATH.mem[INST_ADDR + 8] = {IMM2[11:0], 5'd1, `FNC_LHU, 5'd10, `OPC_LOAD};
    //LHU x10, 2[x1] => x10 = mem[x1 + 0x002] = 32'h0000_face
    `IMEM_PATH.mem[INST_ADDR + 9] = {IMM0[11:0], 5'd1, `FNC_LBU, 5'd11, `OPC_LOAD};
    //LBU x11, 0[x1] => x11 = mem[x1 + 0x000] = 32'h0000_00fe
    `IMEM_PATH.mem[INST_ADDR + 10] = {IMM1[11:0], 5'd1, `FNC_LBU, 5'd12, `OPC_LOAD};
    //LBU x12, 1[x1] => x12 = mem[x1 + 0x001] = 32'h0000_00ca
    `IMEM_PATH.mem[INST_ADDR + 11] = {IMM2[11:0], 5'd1, `FNC_LBU, 5'd13, `OPC_LOAD};
    //LBU x13, 2[x1] => x13 = mem[x1 + 0x002] = 32'h0000_00ce
    `IMEM_PATH.mem[INST_ADDR + 12] = {IMM3[11:0], 5'd1, `FNC_LBU, 5'd14, `OPC_LOAD};
    //LBU x14, 3[x1] => x14 = mem[x1 + 0x003] = 32'h0000_00fa

    `DMEM_PATH.mem[DATA_ADDR] = 32'hface_cafe;

    reset_cpu();

    check_result_rf(5'd2,  32'hface_cafe, "I-Type LW");
    
    check_result_rf(5'd3,  32'hffff_cafe, "I-Type LH 0");
    check_result_rf(5'd4,  32'hffff_face, "I-Type LH 2");

    check_result_rf(5'd5,  32'hffff_fffe, "I-Type LB 0");
    check_result_rf(5'd6,  32'hffff_ffca, "I-Type LB 1");
    check_result_rf(5'd7,  32'hffff_ffce, "I-Type LB 2");
    check_result_rf(5'd8,  32'hffff_fffa, "I-Type LB 3");

    check_result_rf(5'd9, 32'h0000cafe, "I-Type LHU 0");
    check_result_rf(5'd10, 32'h0000face, "I-Type LHU 2");

    check_result_rf(5'd11, 32'h000000fe, "I-Type LBU 0");
    check_result_rf(5'd12, 32'h000000ca, "I-Type LBU 1");
    check_result_rf(5'd13, 32'h000000ce, "I-Type LBU 2");
    check_result_rf(5'd14, 32'h000000fa, "I-Type LBU 3");
end


if (1) begin
    // Test S-Type Insts --------------------------------------------------
    // - SW, SH, SB

    reset();

    `RF_PATH.mem[1]  = 32'hfeed_beef;     //x1
    `RF_PATH.mem[2]  = 32'h3000_0010;  //x2
    `RF_PATH.mem[3]  = 32'h3000_0020;  //x3
    `RF_PATH.mem[4]  = 32'h3000_0030;  //x4
    `RF_PATH.mem[5]  = 32'h3000_0040;  //x5
    `RF_PATH.mem[6]  = 32'h3000_0050;  //x6
    `RF_PATH.mem[7]  = 32'h3000_0060;  //x7
    `RF_PATH.mem[8]  = 32'h3000_0070;  //x8
    `RF_PATH.mem[9]  = 32'h3000_0080;  //x9
    `RF_PATH.mem[10] = 32'h3000_0090; //x10

    IMM0 = 32'h0000_0104;  //Last addr [1:0]
    IMM1 = 32'h0000_0105;
    IMM2 = 32'h0000_0106;
    IMM3 = 32'h0000_0107;
    INST_ADDR = 14'h0000;

    DATA_ADDR0 = (`RF_PATH.mem[2]  + IMM0[11:0]) >> 2;

    DATA_ADDR1 = (`RF_PATH.mem[3]  + IMM0[11:0]) >> 2;
    DATA_ADDR2 = (`RF_PATH.mem[4]  + IMM1[11:0]) >> 2;
    DATA_ADDR3 = (`RF_PATH.mem[5]  + IMM2[11:0]) >> 2;
    DATA_ADDR4 = (`RF_PATH.mem[6]  + IMM3[11:0]) >> 2;

    DATA_ADDR5 = (`RF_PATH.mem[7]  + IMM0[11:0]) >> 2;
    DATA_ADDR6 = (`RF_PATH.mem[8]  + IMM1[11:0]) >> 2;
    DATA_ADDR7 = (`RF_PATH.mem[9]  + IMM2[11:0]) >> 2;
    DATA_ADDR8 = (`RF_PATH.mem[10] + IMM3[11:0]) >> 2;

    `IMEM_PATH.mem[INST_ADDR + 0] = {IMM0[11:5], 5'd1, 5'd2,  `FNC_SW, IMM0[4:0], `OPC_STORE};
    //SW x1, 0x104(x2) => Mem[x2+0x104] = x1 = 0xfeed_beef
    `IMEM_PATH.mem[INST_ADDR + 1] = {IMM0[11:5], 5'd1, 5'd3,  `FNC_SH, IMM0[4:0], `OPC_STORE};
    //SH x1, 0x104(x3) => Mem[x3+0x104] = {16'b0,x1[15:0]} = 0x0000_beef
    `IMEM_PATH.mem[INST_ADDR + 2] = {IMM2[11:5], 5'd1, 5'd5,  `FNC_SH, IMM2[4:0], `OPC_STORE};
    //SH x1, 0x106(x5) => Mem[x5+0x106] = {x1[15:0],16'b0}  = 0xbeef_0000

    `IMEM_PATH.mem[INST_ADDR + 3] = {IMM0[11:5], 5'd1, 5'd7,  `FNC_SB, IMM0[4:0], `OPC_STORE};
    //SB x1, 0x104(x7) => Mem[x7+0x104] = {24'b0,x1[7:0]}  = 0x0000_00ef
    `IMEM_PATH.mem[INST_ADDR + 4] = {IMM1[11:5], 5'd1, 5'd8,  `FNC_SB, IMM1[4:0], `OPC_STORE};
    //SB x1, 0x105(x8) => Mem[x8+0x105] = {16'b0,x1[7:0],8'b0}  = 0x0000_ef00
    `IMEM_PATH.mem[INST_ADDR + 5] = {IMM2[11:5], 5'd1, 5'd9,  `FNC_SB, IMM2[4:0], `OPC_STORE};
    //SB x1, 0x106(x9) => Mem[x9+0x106] = {8'b0,x1[7:0],16'b0}  = 0x00ef_0000
    `IMEM_PATH.mem[INST_ADDR + 6] = {IMM3[11:5], 5'd1, 5'd10, `FNC_SB, IMM3[4:0], `OPC_STORE};
    //SB x1, 0x107(x10) => Mem[x10+0x107] = {x1[7:0],24'b0} = 0xef00_0000

    `DMEM_PATH.mem[DATA_ADDR0] = 0;
    `DMEM_PATH.mem[DATA_ADDR1] = 0;
    `DMEM_PATH.mem[DATA_ADDR3] = 0;
    `DMEM_PATH.mem[DATA_ADDR4] = 0;
    `DMEM_PATH.mem[DATA_ADDR5] = 0;
    `DMEM_PATH.mem[DATA_ADDR6] = 0;
    `DMEM_PATH.mem[DATA_ADDR7] = 0;
    `DMEM_PATH.mem[DATA_ADDR8] = 0;

    reset_cpu();

    check_result_dmem(DATA_ADDR0, 32'hfeed_beef, "S-Type SW");

    check_result_dmem(DATA_ADDR1, 32'h0000_beef, "S-Type SH 1");
    check_result_dmem(DATA_ADDR3, 32'hbeef_0000, "S-Type SH 3");

    check_result_dmem(DATA_ADDR5, 32'h0000_00ef, "S-Type SB 1");
    check_result_dmem(DATA_ADDR6, 32'h0000_ef00, "S-Type SB 2");
    check_result_dmem(DATA_ADDR7, 32'h00ef_0000, "S-Type SB 3");
    check_result_dmem(DATA_ADDR8, 32'hef00_0000, "S-Type SB 4");
end

if (1) begin
    // Test U-Type Insts --------------------------------------------------
    // - LUI, AUIPC
    reset();

    IMM = 32'h9876_abcd;
    INST_ADDR = 14'h0000;
    //RESET_PC = 32'h1000_0000;

    `IMEM_PATH.mem[INST_ADDR + 0] = {IMM[31:12], 5'd7, `OPC_LUI};
    //Current PC = 32'h1000_0000; Next PC = 32'h1000_0004;
    //LUI x7, 0x9876_a_000 => x7 = 0x9876_a000
    `IMEM_PATH.mem[INST_ADDR + 1] = {IMM[31:12], 5'd8, `OPC_AUIPC};
    //Current PC = 32'h1000_0004; Next PC = 32'h1000_0008;
    //AUIPC x8, 0x9876_a_000 => x8 = 0x9876_a000 + PC(0x1000_0004) = 0xa876_a004

    reset_cpu();

    check_result_rf(5'd7,  32'h9876_a000, "U-Type LUI");
    check_result_rf(5'd8,  32'ha876_a004, "U-Type AUIPC");
end

if (1) begin
    // Test J-Type Insts --------------------------------------------------
    // - JAL
    reset();
    //RESET_PC = 32'h1000_0000;

    `RF_PATH.mem[1] = 50;   //x1 = 50
    `RF_PATH.mem[2] = 100; //x2 = 100
    `RF_PATH.mem[3] = 200; //x3 = 200
    `RF_PATH.mem[4] = 300; //x4 = 300

    IMM       = 32'h0000_0aa0; // {IMM[20:1],1'b0} = 0x0aa0
    INST_ADDR = 14'h0000;
    JUMP_ADDR = (32'h1000_0000 + {IMM[20:1], 1'b0}) >> 2;

    `IMEM_PATH.mem[INST_ADDR + 0]   = {IMM[20], IMM[10:1], IMM[11], IMM[19:12], 5'd5, `OPC_JAL};
    //Current PC = 32'h1000_0000; Next PC = 32'h1000_0004;
    //JAL x5, imm[20:1] => PC = PC(0x1000_0000) + {IMM[20:1],1'b0} = 0x1000_0aa0
    //      x5 = Next PC = 0x1000_0004
    `IMEM_PATH.mem[INST_ADDR + 1]   = {`FNC7_0, 5'd2, 5'd1, `FNC_ADD_SUB, 5'd6, `OPC_ARI_RTYPE};
    //Current PC = 32'h1000_0aa0; Next PC = 32'h1000_0aa4; 
    //ADD x6, x1, x2 => x6 = x1 + x2 = 50 + 100 = 150
    //But PC is changed, x6 = 0
    `IMEM_PATH.mem[JUMP_ADDR[13:0]] = {`FNC7_0, 5'd4, 5'd3, `FNC_ADD_SUB, 5'd7, `OPC_ARI_RTYPE};
    //Current PC = 32'h1000_0aa0; Next PC = 32'h1000_0aa4; 
    //ADD x7, x3, x4 => x7 = x3 + x4 = 200 + 300 = 500
    `IMEM_PATH.mem[JUMP_ADDR[13:0] + 1]   = {`FNC7_0, 5'd3, 5'd2, `FNC_ADD_SUB, 5'd8, `OPC_ARI_RTYPE};
    //Current PC = 32'h1000_0aa4; Next PC = 32'h1000_0aa8; 
    //ADD x8, x2, x3 => x8 = x2 + x3 = 100 + 200 = 300

    reset_cpu();

    check_result_rf(5'd5, 32'h1000_0004, "J-Type JAL");
    check_result_rf(5'd7, 500, "J-Type JAL");
    check_result_rf(5'd6, 0, "J-Type JAL");
    check_result_rf(5'd8, 300, "J-Type JAL");
end

if (1) begin
    // Test I-Type JALR Insts ---------------------------------------------
    reset();
    //RESET_PC = 32'h1000_0000;
    `RF_PATH.mem[1] = 32'h1000_0100; //x1
    `RF_PATH.mem[2] = 100;                     //x2 = 100
    `RF_PATH.mem[3] = 300;                     //x3 = 300
    `RF_PATH.mem[4] = 500;                     //x4 = 500

    IMM       = 32'hFFFF_fff0;
    INST_ADDR = 14'h0000;
    JUMP_ADDR = (`RF_PATH.mem[1] + IMM) >> 2;

    `IMEM_PATH.mem[INST_ADDR + 0]   = {IMM[11:0], 5'd1, 3'b000, 5'd5, `OPC_JALR};
    //Current PC = 32'h1000_0000; Next PC = 32'h1000_0004;
    //JALR x5, x1, 0xff0 => PC = x1(0x1000_0100) + 0xff0 = 0x1000_10f0
    //      x5 = Next PC = 0x1000_0004
    `IMEM_PATH.mem[INST_ADDR + 1]   = {`FNC7_0,   5'd2, 5'd4, `FNC_ADD_SUB, 5'd6, `OPC_ARI_RTYPE};
    //Current PC = 32'h1000_10f0; Next PC = 32'h1000_10f4; 
    //ADD x6, x4, x2 => x6 = x4 + x2 = 500 + 100 = 600
    //But PC is changed, x6 = 0
    `IMEM_PATH.mem[JUMP_ADDR[13:0]] = {`FNC7_0,   5'd4, 5'd3, `FNC_ADD_SUB, 5'd7, `OPC_ARI_RTYPE};
    //Current PC = 32'h1000_10f0; Next PC = 32'h1000_10f4; 
    //ADD x7, x3, x4 => x7 = x3 + x4 = 300 + 500 = 800
    `IMEM_PATH.mem[JUMP_ADDR[13:0] + 1]   = {`FNC7_0, 5'd3, 5'd2, `FNC_ADD_SUB, 5'd8, `OPC_ARI_RTYPE};
    //Current PC = 32'h1000_10f4; Next PC = 32'h1000_10f8; 
    //ADD x8, x2, x3 => x8 = x2 + x3 = 100 + 300 = 400

    reset_cpu();

    check_result_rf(5'd5, 32'h1000_0004, "J-Type JALR");
    check_result_rf(5'd7, 800, "J-Type JALR");
    check_result_rf(5'd6, 0, "J-Type JALR");
    check_result_rf(5'd8, 400, "J-Type JALR");
end

if (1) begin
    // Test B-Type Insts --------------------------------------------------
    // - BEQ, BNE, BLT, BGE, BLTU, BGEU

    IMM       = 32'h0000_0FF0;
    INST_ADDR = 14'h0000;
    JUMP_ADDR = (32'h1000_0000 + IMM[12:0]) >> 2;

    BR_TYPE[0]     = `FNC_BEQ;
    BR_NAME_TK1[0] = "B-Type BEQ Taken 1";
    BR_NAME_TK2[0] = "B-Type BEQ Taken 2";
    BR_NAME_NTK[0] = "B-Type BEQ Not Taken";

    //NZCV flag update, RegWrite nop
    BR_TAKEN_OP1[0]  = 300; BR_TAKEN_OP2[0]  = 300;
    //BEQ  IMM  300 - 300 = 0     true,   Btaken = 1
    BR_NTAKEN_OP1[0] = 300; BR_NTAKEN_OP2[0] = 200;
    //BEQ  IMM   300 - 200 = 0    false,   Btaken = 0

    BR_TYPE[1]       = `FNC_BNE;
    BR_NAME_TK1[1]   = "B-Type BNE Taken 1";
    BR_NAME_TK2[1]   = "B-Type BNE Taken 2";
    BR_NAME_NTK[1]   = "B-Type BNE Not Taken";
    //NZCV flag update, RegWrite nop
    BR_TAKEN_OP1[1]  = 300; BR_TAKEN_OP2[1]  = 200;
    //BNE  IMM  300 - 200 != 0     true,   Btaken = 1
    BR_NTAKEN_OP1[1] = 700; BR_NTAKEN_OP2[1] = 700;
    //BNE  IMM   700 - 700 != 0    false,   Btaken = 0

    BR_TYPE[2]       = `FNC_BLT;
    BR_NAME_TK1[2]   = "B-Type BLT Taken 1";
    BR_NAME_TK2[2]   = "B-Type BLT Taken 2";
    BR_NAME_NTK[2]   = "B-Type BLT Not Taken";
    //NZCV flag update, RegWrite nop
    BR_TAKEN_OP1[2]  = 500; BR_TAKEN_OP2[2]  = 700;
    //BLT  IMM  500 - 700 < 0     true,   Btaken = 1
    BR_NTAKEN_OP1[2] = 700; BR_NTAKEN_OP2[2] = 500;
    //BLT  IMM   300 - 200 < 0    false,   Btaken = 0

    BR_TYPE[3]       = `FNC_BGE;
    BR_NAME_TK1[3]   = "B-Type BGE Taken 1";
    BR_NAME_TK2[3]   = "B-Type BGE Taken 2";
    BR_NAME_NTK[3]   = "B-Type BGE Not Taken";
    //NZCV flag update, RegWrite nop
    BR_TAKEN_OP1[3]  = 800; BR_TAKEN_OP2[3]  = 300;
    //BGE  IMM  800 - 300 >= 0     true,   Btaken = 1
    BR_NTAKEN_OP1[3] = 300; BR_NTAKEN_OP2[3] = 800;
    //BGE  IMM   300 - 800 >= 0    false,   Btaken = 0

    BR_TYPE[4]       = `FNC_BLTU;
    BR_NAME_TK1[4]   = "B-Type BLTU Taken 1";
    BR_NAME_TK2[4]   = "B-Type BLTU Taken 2";
    BR_NAME_NTK[4]   = "B-Type BLTU Not Taken";
    //NZCV flag update, RegWrite nop
    BR_TAKEN_OP1[4]  = 32'h0000_000a; BR_TAKEN_OP2[4]  = 32'haaaa_0000;
    //BLTU IMM 0x0000_0001 - 0xaaaa_0000 < 0 true, Btaken = 1 unsigned
    BR_NTAKEN_OP1[4] = 32'haaaa_0000; BR_NTAKEN_OP2[4] = 32'h0000_000a;
    //BLTU IMM 0xaaaa_0000 - 0x0000_0001 < 0 false, Btaken = 0 unsigned

    BR_TYPE[5]       = `FNC_BGEU;
    BR_NAME_TK1[5]   = "B-Type BGEU Taken 1";
    BR_NAME_TK2[5]   = "B-Type BGEU Taken 2";
    BR_NAME_NTK[5]   = "B-Type BGEU Not Taken";
    //NZCV flag update, RegWrite nop
    BR_TAKEN_OP1[5]  = 32'haaaa_0000; BR_TAKEN_OP2[5]  = 32'h0000_000a;
    //BGEU IMM 0x0000_0001 - 0xaaaa_0000 < 0 true, Btaken = 1 unsigned
    BR_NTAKEN_OP1[5] = 32'h0000_000a; BR_NTAKEN_OP2[5] = 32'haaaa_0000;
    //BGEU IMM 0xaaaa_0000 - 0x0000_0001 < 0 false, Btaken = 0 unsigned
    for (i = 0; i < 6; i = i + 1) begin
      reset();

      `RF_PATH.mem[1] = BR_TAKEN_OP1[i];
      `RF_PATH.mem[2] = BR_TAKEN_OP2[i];
      `RF_PATH.mem[3] = 70;
      `RF_PATH.mem[4] = 707;
      `RF_PATH.mem[9] = 7;
/*
    `IMEM_PATH.mem[INST_ADDR + 0]   = {IMM[11:0], 5'd1, 3'b000, 5'd5, `OPC_JALR};
    //Current PC = 32'h1000_0000; Next PC = 32'h1000_0004;
    //JALR x5, x1, 0xff0 => PC = x1(0x1000_0100) + 0xff0 = 0x1000_10f0
    //      x5 = Next PC = 0x1000_0004
    `IMEM_PATH.mem[INST_ADDR + 1]   = {`FNC7_0,   5'd2, 5'd4, `FNC_ADD_SUB, 5'd6, `OPC_ARI_RTYPE};
    //Current PC = 32'h1000_10f0; Next PC = 32'h1000_10f4; 
    //ADD x6, x4, x2 => x6 = x4 + x2 = 500 + 100 = 600
    //But PC is changed, x6 = 0
    `IMEM_PATH.mem[JUMP_ADDR[13:0]] = {`FNC7_0,   5'd4, 5'd3, `FNC_ADD_SUB, 5'd7, `OPC_ARI_RTYPE};
    //Current PC = 32'h1000_10f0; Next PC = 32'h1000_10f4; 
    //ADD x7, x3, x4 => x7 = x3 + x4 = 300 + 500 = 800
    `IMEM_PATH.mem[JUMP_ADDR[13:0] + 1]   = {`FNC7_0, 5'd3, 5'd2, `FNC_ADD_SUB, 5'd8, `OPC_ARI_RTYPE};
    //Current PC = 32'h1000_10f4; Next PC = 32'h1000_10f8; 
    //ADD x8, x2, x3 => x8 = x2 + x3 = 100 + 300 = 400
*/


      // Test branch taken
      `IMEM_PATH.mem[INST_ADDR + 0]   = {IMM[12], IMM[10:5], 5'd2, 5'd1, BR_TYPE[i], IMM[4:1], IMM[11], `OPC_BRANCH};
      //Current PC = 32'h1000_0000; Next PC = 32'h1000_0004;
      //B  x1, x2 if true, Branch  PC = PC + 0xff0
      `IMEM_PATH.mem[INST_ADDR + 1]   = {`FNC7_0, 5'd4, 5'd3, `FNC_ADD_SUB, 5'd5, `OPC_ARI_RTYPE};
      //Current PC = 32'h1000_0ff0; Next PC = 32'h1000_0ff4;
      //ADD x5, x3, x4 => x5 = x3 + x4 = 70 + 707 = 777
      //But PC is changed, x5 = 0
      `IMEM_PATH.mem[JUMP_ADDR[13:0]] = {`FNC7_0, 5'd4, 5'd3, `FNC_ADD_SUB, 5'd6, `OPC_ARI_RTYPE};
      //Current PC = 32'h1000_0ff0; Next PC = 32'h1000_0ff4;
      //ADD x6, x3, x4 => x6 = x3 + x4 = 70 + 707 = 777
      `IMEM_PATH.mem[JUMP_ADDR[13:0] + 1] = {`FNC7_0, 5'd9, 5'd3, `FNC_ADD_SUB, 5'd7, `OPC_ARI_RTYPE};
      //Current PC = 32'h1000_0ff4; Next PC = 32'h1000_0ff8;
      //ADD x7, x3, x9 => x7 = x3 + x9 = 70 + 7 = 77

      reset_cpu();

      check_result_rf(5'd5, 0,   BR_NAME_TK1[i]);
      check_result_rf(5'd6, 777, BR_NAME_TK2[i]);
      check_result_rf(5'd7, 77, BR_NAME_TK2[i]);

      reset();

      `RF_PATH.mem[1] = BR_NTAKEN_OP1[i];
      `RF_PATH.mem[2] = BR_NTAKEN_OP2[i];
      `RF_PATH.mem[3] = 70;
      `RF_PATH.mem[4] = 707;

      // Test branch not taken
      `IMEM_PATH.mem[INST_ADDR + 0] = {IMM[12], IMM[10:5], 5'd2, 5'd1, BR_TYPE[i], IMM[4:1], IMM[11], `OPC_BRANCH};
      //Current PC = 32'h1000_0000; Next PC = 32'h1000_0004;
      //B  x1, x2 if false,  PC = Next PC
      `IMEM_PATH.mem[INST_ADDR + 1] = {`FNC7_0, 5'd4, 5'd3, `FNC_ADD_SUB, 5'd5, `OPC_ARI_RTYPE};
      //Current PC = 32'h1000_0004; Next PC = 32'h1000_0008;
      //ADD x5, x3, x4 => x5 = x3 + x4 = 70 + 707 = 777

      reset_cpu();
      check_result_rf(5'd5, 777, BR_NAME_NTK[i]);
    end
end


    // ... what else?
    all_tests_passed = 1'b1;

    repeat (100) @(posedge clk);
    $display("All tests passed!");
    $finish();
  end

endmodule
