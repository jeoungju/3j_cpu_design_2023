module p_d_DE(
    port_list
);
    
endmodule